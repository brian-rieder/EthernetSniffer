// File name:   comparator.sv
// Updated:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: comparator

module comparator
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
