// File name:   controller.sv
// Updated:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: controller

module controller
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
