// File name:   avalon_slave_controller.sv
// Created:     05 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: avalon_slave_controller

module avalon_slave_controller
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
