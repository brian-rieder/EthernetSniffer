// File name:   result_address_fsm.sv
// Created:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: result_address_fsm

module result_address_fsm
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
