// File name:   result_address_lookup.sv
// Updated:     16 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: result_address_lookup

module result_address_lookup
(
  // port declaration
);

endmodule
