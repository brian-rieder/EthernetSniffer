// File name:   comparator.sv
// Created:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: comparator

module comparator
#(
  // parameter declaration
)
(
  // port declaration
  input wire [31:0]data
  output wire [31:0]data
);

endmodule
