// File name:   tmp.sv
// Created:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: tmp

module tmp
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
