// File name:   comparator_addresses.sv
// Created:     04 November 2015
// Authors:     Brian Rieder 
//              Catie Cowden 
//              Shaughan Gladden
// Description: comparator_addresses

module comparator_addresses
#(
  // parameter declaration
)
(
  // port declaration
);

endmodule
